module CPU_WrapperV2 (
    input clk,
    input rstn,
    input [7 : 0] I_Port,
    input [7 : 0] I_Port,
    output [7 : 0] O_Port
);



endmodule