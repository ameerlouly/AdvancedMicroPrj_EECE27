module CPU_Wrapper1(
    input
    output
);

endmodule